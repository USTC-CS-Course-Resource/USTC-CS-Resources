module test(	//ģ������
    input in,	//�����ź�����
    output out,	//����ź�����
    output out_n);
    //���ڴ������ڲ�����
    /*******����Ϊ�߼���������******/
    assign out = in;
    assign out_n = ~in;
    /*******�߼��������ֽ���******/
endmodule   //ģ���������ؼ���

